module qam_64 #(
    parameter INPUT_DATA_WIDTH = 12,                     // Width of the input data
    parameter OUTPUT_DATA_WIDTH_I = 16,                  // Width of the I channel output data
    parameter OUTPUT_DATA_WIDTH_Q = 16,                  // Width of the Q channel output data
    parameter QAM64_AMPLITUDE = 16'b0001001111000000    // Amplitude of the QAM-64 signal
) (
    input clk,                                          // Clock input
    input enable,                                       // Enable signal to activate modulation
    input [INPUT_DATA_WIDTH-1:0] data_in,               // Input data to be modulated
    output reg signed [OUTPUT_DATA_WIDTH_I-1:0] channel_i [0:(INPUT_DATA_WIDTH/6)-1],  // Output I channel
    output reg signed [OUTPUT_DATA_WIDTH_Q-1:0] channel_q [0:(INPUT_DATA_WIDTH/6)-1]   // Output Q channel
);

    integer i;  // Declare loop counter

    always @(*) begin
        // Loop through each symbol of the input data (6 bits per symbol for QAM-64)
        for (i = 0; i < (INPUT_DATA_WIDTH / 6); i = i + 1) begin
            // Calculate in-phase (I) channel using QAM-64 modulation formula
            // QAM64_AMPLITUDE * (1 - 2 * data_in[6*i]) * (4 - (1 - 2 * data_in[6*i + 2]) * (2 - (1 - 2 * data_in[6*i + 4])))
            channel_i[i] = enable ? QAM64_AMPLITUDE * (1 - 2 * data_in[6*i]) * (4 - (1 - 2 * data_in[6*i + 2]) * (2 - (1 - 2 * data_in[6*i + 4]))) : 'd0;
            
            // Calculate quadrature (Q) channel using QAM-64 modulation formula
            // QAM64_AMPLITUDE * (1 - 2 * data_in[6*i + 1]) * (4 - (1 - 2 * data_in[6*i + 3]) * (2 - (1 - 2 * data_in[6*i + 5])))
            channel_q[i] = enable ? QAM64_AMPLITUDE * (1 - 2 * data_in[6*i + 1]) * (4 - (1 - 2 * data_in[6*i + 3]) * (2 - (1 - 2 * data_in[6*i + 5]))) : 'd0;
        end
    end
    
endmodule
